LIBRARY ieee;
USE ieee.std_logic_1164.all;

--Simple module that connects the SW switches to the LEDR lights

ENTITY part1 IS
	PORT(SW		:IN 		STD_LOGIC_VECTOR(9 DOWNTO 0);
		  LEDR	:OUT		STD_LOGIC_VECTOR(9 DOWNTO 0));
END part1;

ARCHITECTURE Behaviour OF part1 IS
BEGIN
	LEDR <= SW;
END Behaviour;
		  
		  